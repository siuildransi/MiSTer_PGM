module top (
    input         FPGA_CLK1_50,
    input         FPGA_CLK2_50,
    input         FPGA_CLK3_50,

    inout  [35:0] GPIO,
    inout  [14:0] HPS_DDR3_ADDR,
    inout  [2:0]  HPS_DDR3_BA,
    inout         HPS_DDR3_CAS_N,
    inout         HPS_DDR3_CKE,
    inout         HPS_DDR3_CK_N,
    inout         HPS_DDR3_CK_P,
    inout         HPS_DDR3_CS_N,
    inout  [3:0]  HPS_DDR3_DM,
    inout  [31:0] HPS_DDR3_DQ,
    inout  [3:0]  HPS_DDR3_DQS_N,
    inout  [3:0]  HPS_DDR3_DQS_P,
    inout         HPS_DDR3_ODT,
    inout         HPS_DDR3_RAS_N,
    inout         HPS_DDR3_RESET_N,
    inout         HPS_DDR3_RZQ,
    inout         HPS_DDR3_WE_N,

    output [12:0] SDRAM_ADDR,
    output [1:0]  SDRAM_BA,
    output        SDRAM_CAS_N,
    output        SDRAM_CKE,
    output        SDRAM_CLK,
    output        SDRAM_CS_N,
    inout  [15:0] SDRAM_DQ,
    output        SDRAM_LDQM,
    output        SDRAM_RAS_N,
    output        SDRAM_UDQM,
    output        SDRAM_WE_N,

    output        VGA_BLANK_N,
    output [7:0]  VGA_B,
    output        VGA_CLK,
    output [7:0]  VGA_G,
    output        VGA_HS,
    output [7:0]  VGA_R,
    output        VGA_SYNC_N,
    output        VGA_VS
);

// --- Clocks ---
wire clk_20m, clk_8m, clk_sys;
// For now, we'll use simple clock dividers for placeholders
// A proper PLL should be added in sys/pll.qip
reg [1:0] div20;
always @(posedge FPGA_CLK1_50) div20 <= div20 + 2'd1;
assign clk_20m = div20[1]; // ~12.5MHz (placeholder)

reg [2:0] div8;
always @(posedge FPGA_CLK1_50) div8 <= div8 + 3'd1;
assign clk_8m = div8[2];  // ~6.25MHz (placeholder)

assign clk_sys = FPGA_CLK1_50;

// --- Reset ---
wire reset;

// --- Video System ---
wire [7:0] r, g, b;
wire hs, vs, blank_n;

pgm_video video_gen (
    .clk(FPGA_CLK1_50), // 50MHz for standard VGA placeholder
    .reset(reset),
    .hs(hs),
    .vs(vs),
    .r(r),
    .g(g),
    .b(b),
    .blank_n(blank_n)
);

// --- sys_top MiSTer Framework ---
wire ioctl_download, ioctl_wr;
wire [26:0] ioctl_addr;
wire [15:0] ioctl_dout;
wire [7:0]  ioctl_index;

sys_top mister_sys (
    .FPGA_CLK1_50(FPGA_CLK1_50),
    .FPGA_CLK2_50(FPGA_CLK2_50),
    .FPGA_CLK3_50(FPGA_CLK3_50),

    .SDRAM_A(SDRAM_ADDR),
    .SDRAM_DQ(SDRAM_DQ),
    .SDRAM_DQML(SDRAM_LDQM),
    .SDRAM_DQMH(SDRAM_UDQM),
    .SDRAM_nWE(SDRAM_WE_N),
    .SDRAM_nCAS(SDRAM_CAS_N),
    .SDRAM_nRAS(SDRAM_RAS_N),
    .SDRAM_nCS(SDRAM_CS_N),
    .SDRAM_BA(SDRAM_BA),
    .SDRAM_CLK(SDRAM_CLK),
    .SDRAM_CKE(SDRAM_CKE),

    .VGA_R(r[7:2]),
    .VGA_G(g[7:2]),
    .VGA_B(b[7:2]),
    .VGA_HS(hs),
    .VGA_VS(vs),
    .VGA_EN(blank_n),

    // ioctl ROM loading
    .ioctl_download(ioctl_download),
    .ioctl_addr(ioctl_addr),
    .ioctl_dout(ioctl_dout),
    .ioctl_wr(ioctl_wr),
    .ioctl_index(ioctl_index)
);

// --- PGM Core Instance ---
PGM pgm_core (
    .fixed_20m_clk(clk_20m),
    .fixed_8m_clk(clk_8m),
    .reset(reset || ioctl_download), // Reset core during download

    // ioctl
    .ioctl_download(ioctl_download),
    .ioctl_wr(ioctl_wr),
    .ioctl_addr(ioctl_addr),
    .ioctl_dout(ioctl_dout),
    .ioctl_index(ioctl_index),

    // Placeholder connections
    .cpu68k_din(16'hFFFF),
    .cpuz80_din(8'hFF),
    .cpu68k_dtack_n(1'b0)
);

assign reset = ~KEY[0]; // Temporary reset from Button 0

endmodule
